// Code your testbench here
// or browse Examples


`include "uvm_macros.svh"
import uvm_pkg ::*;

module tb;
  initial begin
    `uvm_info("TB_TOP", "Hello World", UVM_NONE);
  end
endmodule

